** sch_path: /foss/designs/libs/tb_single_mos/tb_single_nmos.sch
**.subckt tb_single_nmos
VB net2 GND 0.91
VDD net1 GND 3.3
XM1 net1 GND net2 GND unit_nmos M=1
**** begin user architecture code

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical



.control
    save all
    op
    show all
.endc


**** end user architecture code
**.ends

* expanding   symbol:  libs/core_single_mos/unit_nmos/unit_nmos.sym # of pins=4
** sym_path: /foss/designs/libs/core_single_mos/unit_nmos/unit_nmos.sym
** sch_path: /foss/designs/libs/core_single_mos/unit_nmos/unit_nmos.sch
.subckt unit_nmos drain sub gate source
*.iopin drain
*.iopin source
*.iopin sub
*.iopin gate
XM1 drain gate source sub nfet_03v3 L=0.5u W=12u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m={M}
**** begin user architecture code

.param M=1

**** end user architecture code
.ends

.GLOBAL GND
.end
