** sch_path: /foss/designs/libs/tb_current_mirror/tb_nmos_current_mirror.sch
**.subckt tb_nmos_current_mirror
X_NCM net7 net6 net5 net4 net3 net1 GND nmos_current_mirror
VDD net2 GND 3.3
Ibias net2 net1 100u
VOUT out GND 3.3
Viout1x out net3 0
.save i(viout1x)
Viout2x out net4 0
.save i(viout2x)
Viout4x out net5 0
.save i(viout4x)
Viout16x out net7 0
.save i(viout16x)
Viout8x out net6 0
.save i(viout8x)
**** begin user architecture code

.include /foss/pdks/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /foss/pdks/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical



.control
    save all

    * Operating Point Analysis
    op
    show all > op.log

    * DC Sweep
    dc VOUT 0 3.3 10m
    plot i(viout1x) i(viout2x) i(viout4x) i(viout8x) i(viout16x) vs v(out)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  libs/core_current_mirror/nmos_current_mirror/nmos_current_mirror.sym # of pins=7
** sym_path: /foss/designs/libs/core_current_mirror/nmos_current_mirror/nmos_current_mirror.sym
** sch_path: /foss/designs/libs/core_current_mirror/nmos_current_mirror/nmos_current_mirror.sch
.subckt nmos_current_mirror 16x_I_ref 8x_I_ref 4x_I_ref 2x_I_ref 1x_I_ref I_ref VSS
*.iopin I_ref
*.iopin VSS
*.iopin 1x_I_ref
*.iopin 2x_I_ref
*.iopin 4x_I_ref
*.iopin 8x_I_ref
*.iopin 16x_I_ref
XIREF I_ref VSS I_ref VSS unit_nmos M=1
X1x 1x_I_ref VSS I_ref VSS unit_nmos M=1
X2x 2x_I_ref VSS I_ref VSS unit_nmos M=2
X4x 4x_I_ref VSS I_ref VSS unit_nmos M=4
X8x 8x_I_ref VSS I_ref VSS unit_nmos M=8
X16x 16x_I_ref VSS I_ref VSS unit_nmos M=16
.ends


* expanding   symbol:  libs/core_single_mos/unit_nmos/unit_nmos.sym # of pins=4
** sym_path: /foss/designs/libs/core_single_mos/unit_nmos/unit_nmos.sym
** sch_path: /foss/designs/libs/core_single_mos/unit_nmos/unit_nmos.sch
.subckt unit_nmos drain sub gate source
*.iopin drain
*.iopin source
*.iopin sub
*.iopin gate
XM1 drain gate source sub nfet_03v3 L=0.5u W=12u nf=2 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m={M}
**** begin user architecture code

.param M=1

**** end user architecture code
.ends

.GLOBAL GND
.end
